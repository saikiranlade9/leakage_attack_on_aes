`include "timescale.v"

module master_wrapper_top(PCLK, PRESETn, PADDR, PWDATA, PPROT, PSELx, PENABLE, PWRITE, PSTRB, PREADY, PSLVERR, PRDATA,
                      host_instruction, host_data, start, out, operation_done);

`include "config_pkg.vh"  
   
    //Global Input signals and inputs from host
    input wire  [HOST_INSTRUCT_SIZE-1:0]    host_instruction;
    input wire  [MAX_INPUT_DATA_SIZE-1:0]   host_data;
    input wire                              start;
   
    // Global Clock Signal 
    input   wire    PCLK;
    // Global Reset Signal. This Signal is Active LOW 
    input   wire    PRESETn;
           
    // Write address (generated by master wrapper, acceped by Slave)
    output  wire    [APB_ADDR_WIDTH-1 : 0]  PADDR;
    // Write data (issued by master, acceped by Slave)
    output  wire    [APB_DATA_WIDTH-1 : 0]  PWDATA;
    // This signal indicates the privilege and
    // security level of the transaction
    output  wire    [2 : 0]   PPROT;
    // It indicates that the slave device to be selected
    output  wire    [PSELx_WIDTH-1 :0]   PSELx;
    // Enable. This signal indicates the second and subsequent cycles
    // of an APB transfer
    output  wire    PENABLE;
    // This signal indicates an APB write access when HIGH and an APB 
    // read access when LOW.
    output  wire    PWRITE;
    // It enables sparse data transfer on the write data bus.
    output  wire    [APB_STROBE_WIDTH-1 : 0]   PSTRB;
    
    // Indicates completion of an APB transfer 
    input  wire     PREADY;
    // Indicates a transfer failure 
    input  wire     PSLVERR;
    // Read data (issued by slave)
    input  wire     [APB_DATA_WIDTH-1 : 0]  PRDATA;
    
    //output signals to host
    output wire operation_done;
	output wire [MAX_OUTPUT_DATA_SIZE-1:0] out;
	
	 // This signal, from master,  indicates initiation of a transaction
    wire     init_transaction;
    // AES input text 
    wire    [AES_TEXT_IN_WIDTH-1 : 0] aes_text_in;
    // AES key
    wire    [AES_KEY_WIDTH-1 : 0] aes_key;
    // Input to HASH 
    wire    [HASH_IN_WIDTH-1 : 0] hash_in;
    
    // This signal, from master, indicates the type of transaction master IP
    // wants to perform
    wire   [OPERATION_TYPE_WIDTH-1 : 0]  operation_type;
    
    //outputs to HOST interface 
    //output           input_data_transfer_complete,
    // This signal indicates that the requested data is ready to be read
    wire    data_input_ready;
    // This signal indicates that the provided data is written to respective slave registers
    wire    write_complete;  
    
    // Encrypted data from AES cipher 
    wire    [AES_CIPH_OUT_WIDTH-1 : 0] encrypt_output_data;
    // Decrypted plain text from AES inv cipher
    wire    [AES_INV_CIPH_OUT_WIDTH-1 : 0] decrypt_output_data;
    // Output from HASH
    wire    [HASH_OUT_WIDTH-1 :0] hash_output;

    // This signal, from slave IP, indicates that the transaction failed
    wire    txn_error;
    
    // Operating states for the APB FSM
    reg [1:0] state, next_state;
    
    reg [1:0] aes_encrypt_write_state;
    reg [1:0] aes_encrypt_read_state;
    reg [2:0] aes_decrypt_write_state;
    reg [1:0] aes_decrypt_read_state;
    reg [1:0] hash_write_state;
    reg [1:0] hash_read_state;
    
    // APB4 signals 
    reg [APB_ADDR_WIDTH-1 : 0]  paddr_r, paddr;
    reg [2 : 0]                     pselx_r, pselx;
    reg                             pwrite_r, pwrite;
    reg [APB_DATA_WIDTH-1 : 0]  pwdata_r, pwdata;
    reg                             pstrb_r, pstrb;
    reg                             pprot_r, pprot;
    reg                             penable;
    
    // signals for Wrapper FSM
    reg         en_transfer_r;
    reg [4:0]   count;
    reg [PSELx_WIDTH-1:0]   slave_sel;
    wire        en_transfer;
    reg         operation_complete_r;
    
    reg         delay_reg0, delay_reg1, delay_reg2, delay_reg3;  
    // registers to store the outputs from each slave
    reg                                 write_complete_r;
    reg                                 data_input_ready_r;
    
    // registers to sample inputs from respective slaves upon completion of a transaction.
    reg [AES_CIPH_OUT_WIDTH-1 : 0]      encrypt_output_data_r;
    reg [AES_INV_CIPH_OUT_WIDTH-1 : 0]  decrypt_output_data_r;
    reg [HASH_OUT_WIDTH-1 : 0]          hash_output_r;
    
    // registers to sample inputs from the master upon initiation of a transaction.
    reg [AES_KEY_WIDTH-1 : 0]       aes_key_r;
    reg [AES_TEXT_IN_WIDTH-1 : 0]   aes_text_in_r;
    reg [HASH_IN_WIDTH-1 : 0]       hash_in_r;
 
    
    
    localparam reg [3:0]    AES_ENCRYPT_WRITE = 5'h01,
                            AES_ENCRYPT_READ = 5'h09,
                            AES_DECRYPT_WRITE = 5'h02,
                            AES_DECRYPT_READ= 5'h0a,
                            HASH_WRITE = 5'h05,
                            HASH_READ = 5'h0d;

    
    localparam reg [1:0]    INIT = 2'b00,
                            IDLE = 2'b01,
                            SETUP = 2'b10,
                            ACCESS = 2'b11;
                            
    localparam reg [1:0]    WRITE_AES_ENCRYPT_INIT = 2'b00,
                            WRITE_AES_ENCRYPT_KEY = 2'b01,
                            WRITE_AES_ENCRYPT_DATA_IN = 2'b10,
                            WRITE_AES_ENCRYPT_LOAD = 2'b11;
                            
    localparam reg [1:0]    READ_AES_ENCRYPT_INIT = 2'b00,
                            READ_AES_ENCRYPT_DATA = 2'b01,
                            READ_AES_ENCRYPT_DONE = 2'b10;
                            
    localparam reg [2:0]    WRITE_AES_DECRYPT_INIT = 3'b000,
                            WRITE_AES_DECRYPT_KEY = 3'b001,
                            WRITE_AES_DECRYPT_DATA_IN = 3'b010,
                            WRITE_AES_DECRYPT_LOAD = 3'b011,
                            WRITE_AES_DECRYPT_K_LOAD = 3'b100;
 
    localparam reg [1:0]    READ_AES_DECRYPT_INIT = 2'b00,
                            READ_AES_DECRYPT_DATA = 2'b01,
                            READ_AES_DECRYPT_DONE = 2'b10;
                            
    localparam reg [1:0]    WRITE_HASH_INIT = 2'b00,
                            WRITE_HASH_DATA_IN = 2'b01,
                            WRITE_HASH_GO = 2'b10; 
                            
    localparam reg [1:0]    READ_HASH_INIT = 2'b00,
                            READ_HASH_DATA = 2'b01,
                            READ_HASH_DONE = 2'b10;    
       
    assign en_transfer = en_transfer_r;
    
    assign encrypt_output_data = encrypt_output_data_r;
    assign decrypt_output_data = decrypt_output_data_r;
    assign hash_output = hash_output_r;
    
       
    assign data_input_ready = data_input_ready_r;
    assign write_complete = write_complete_r;
    assign PADDR = paddr;
    assign PSELx = pselx;
    assign PWRITE = pwrite;
    assign PWDATA = pwdata;
    assign PSTRB = pstrb;
    assign PPROT = pprot;
    assign PENABLE = penable;               
    
    assign txn_error = PREADY ? PSLVERR : 0;
 
    // counter to keep track of transactions and generate addresses.                
    always@(posedge PCLK or negedge PRESETn)
    begin
        if(PRESETn == 1'b0)
            count <= 0;
        else
        begin
            if( (operation_complete_r == 1'b1) | (init_transaction == 1'b0))
                count <= 0;
            else if( (state == SETUP) && (en_transfer == 1'b1))
            begin
                count <= count + 5'h01;
            end
        end
    end
    
    always@(posedge PCLK or negedge PRESETn)
    begin
        if(PRESETn == 1'b0)
        begin
            delay_reg0 <= 0;
            delay_reg1 <= 0;
            delay_reg2 <= 0;
            delay_reg3 <= 0;
        end
        else if(init_transaction == 1'b1)
        begin
            delay_reg0 <= 1;
            delay_reg1 <= delay_reg0;
            delay_reg2 <= delay_reg1;
            delay_reg3 <= delay_reg2;
        end
        else
        begin
            delay_reg0 <= 0;
            delay_reg1 <= 0;
            delay_reg2 <= 0;
            delay_reg3 <= 0;
        end 
    end
    

    // assign appropriate value to slave sel based on the type of operation requested
    always@(*)
    begin
        case(operation_type)
            AES_ENCRYPT_WRITE:  slave_sel = 3'b001;
            AES_ENCRYPT_READ:   slave_sel = 3'b001;
            AES_DECRYPT_WRITE:  slave_sel = 3'b001;
            AES_DECRYPT_READ:   slave_sel = 3'b001;
            HASH_WRITE:         slave_sel = 3'b010;
            HASH_READ:          slave_sel = 3'b010;
            default:            slave_sel = 3'b000;
        endcase
    end

    // Wrapper FSMD
    always@(posedge PCLK or negedge PRESETn)
    begin
        if( PRESETn == 1'b0 )
            begin
                paddr_r <= 0;
                pprot_r <= 0;
                pselx_r <= 0;
                pwrite_r <= 0;
                pwdata_r <= 0;
                pstrb_r <= 0;
                
                en_transfer_r <= 0;
                operation_complete_r <= 0;
                write_complete_r <= 0;
                data_input_ready_r <= 0;
                
                aes_encrypt_write_state <= 0;
                aes_encrypt_read_state <= 0;
                aes_decrypt_write_state <= 0;
                aes_decrypt_read_state <= 0;
                hash_write_state <= 0;
                hash_read_state <= 0;
                
                encrypt_output_data_r <= 0;
                decrypt_output_data_r <= 0;
                hash_output_r <= 0;
                
                aes_key_r <= 0;
                aes_text_in_r <= 0;
                hash_in_r <= 0;
            end
            
        
        else if( init_transaction == 1'b1 )
            begin
                //control signals generated will be HIGH only for one cycle
                write_complete_r <= 0;
                data_input_ready_r <= 0;
                operation_complete_r <= 0;
                case(operation_type)

 //#################################### AES ENCRYPT #################################################                    
                    AES_ENCRYPT_WRITE:
                        begin
                            pselx_r <= slave_sel;
                            pwrite_r <= 1'b1;
                            case(aes_encrypt_write_state)
                                
                                WRITE_AES_ENCRYPT_INIT:
                                begin
                                    aes_key_r <= AES_KEY;
                                    aes_text_in_r <= aes_text_in;
                                    if( (PREADY == 1'b1) && (slave_sel != 0) && (write_complete != 1) )
                                        aes_encrypt_write_state <= WRITE_AES_ENCRYPT_KEY;
                                      
                                end
                                
                                WRITE_AES_ENCRYPT_KEY:
                                begin
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b00100) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + count*4;
                                            pwdata_r <= aes_key_r[APB_DATA_WIDTH-1 : 0];
                                            if(delay_reg1 == 1)
                                            begin
                                                aes_key_r <= aes_key_r >> APB_DATA_WIDTH;
                                            end
                                            en_transfer_r <= 1;
                                        end 
                                    else if( (count == 5'b00011) && (state == SETUP))
                                        begin
                                            //en_transfer_r <= 1'b0;
                                            aes_encrypt_write_state <= WRITE_AES_ENCRYPT_DATA_IN;                                
                                        end                                                        
                                end
                                
                                WRITE_AES_ENCRYPT_DATA_IN:
                                begin
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b01000) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + count*4;
                                            pwdata_r <= aes_text_in_r[APB_DATA_WIDTH-1 : 0];
                                            aes_text_in_r <= aes_text_in_r >> APB_DATA_WIDTH;
                                            en_transfer_r <= 1'b1;
                                        end 
                                    else if( (count == 5'b00111) && (state == SETUP) )
                                        begin
                                            //en_transfer_r <= 1'b0;
                                            aes_encrypt_write_state <= WRITE_AES_ENCRYPT_LOAD;                                
                                        end                                                        
                                end
                                
                                WRITE_AES_ENCRYPT_LOAD:
                                begin
                                    pstrb_r <= 4'b0000;
                                    
                                    if( (count < 5'b01001) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + count*4;
                                            pwdata_r <= 32'h00000001;
                                            en_transfer_r <= 1'b1;
                                        end 
                                        
                                    else if( (count == 5'b01001) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + (count - 5'h01)*4;
                                            pwdata_r <= 32'h0000_0000;
                                            en_transfer_r <= 1'b1;
                                        end
                                        
                                    else if( (count == 5'b01001) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 1'b0;
                                            //pselx_r <= 0;
                                            operation_complete_r <= 1;
                                        end
                                     
                                    else if( (count == 5'b01001) && (PREADY == 1'b1) )
                                        begin
                                            pselx_r <= 0;
                                        end
                                        
                                    else if( (count == 5'b01010) && (PREADY == 1'b1) )
                                        begin
                                            write_complete_r <= 1;
                                            aes_encrypt_write_state <= WRITE_AES_ENCRYPT_INIT;                                    
                                        end 
                                                                                            
                                end
                                
                                default:
                                begin
                                    aes_encrypt_write_state <= WRITE_AES_ENCRYPT_INIT;
                                end                        
                              
                            endcase   
                        end
                        
                        
                    AES_ENCRYPT_READ:
                        begin
                            case(aes_encrypt_read_state)
                                
                                READ_AES_ENCRYPT_INIT:
                                begin
                                    if( (PREADY == 1) && (slave_sel != 0) )
                                        aes_encrypt_read_state <= READ_AES_ENCRYPT_DATA;
                                    en_transfer_r <= 0;
                                end
                                
                                READ_AES_ENCRYPT_DATA:
                                begin
                                    pselx_r <= slave_sel;
                                    pwrite_r <= 1'b0;
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b00100) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_READ_00 + count*4;
                                            encrypt_output_data_r <= {PRDATA, encrypt_output_data[AES_CIPH_OUT_WIDTH-1 : APB_DATA_WIDTH]};
                                            en_transfer_r <= 1'b1;
                                        end
                                    else if( (count == 5'b00011) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 0;
                                        end
                                        
                                    else if( (count == 5'b00100) && (PREADY == 1'b1) )
                                            begin
                                                encrypt_output_data_r <= {PRDATA, encrypt_output_data[AES_CIPH_OUT_WIDTH-1 : APB_DATA_WIDTH]};
                                                aes_encrypt_read_state <= READ_AES_ENCRYPT_DONE;   
                                            end 
                                end 
                                READ_AES_ENCRYPT_DONE:
                                begin
                                    pselx <= 0;
                                    operation_complete_r <= 1;
                                    data_input_ready_r <= 1;
                                    aes_encrypt_read_state <= READ_AES_ENCRYPT_INIT;
                                end
                            endcase
                        end

 //#################################### AES DECRYPT ################################################# 
                        
                    AES_DECRYPT_WRITE:
                        begin
                            pselx_r <= slave_sel;
                            pwrite_r <= 1'b1;
                            case(aes_decrypt_write_state)
                                
                                WRITE_AES_DECRYPT_INIT:
                                begin
                                    aes_key_r <= AES_KEY;
                                    aes_text_in_r <= aes_text_in;
                                    if( (PREADY == 1'b1) && (slave_sel != 0) && (write_complete != 1) )
                                        aes_decrypt_write_state <= WRITE_AES_DECRYPT_KEY;
                                      
                                end
                                
                                WRITE_AES_DECRYPT_KEY:
                                begin
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b00100) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + count*4;
                                            pwdata_r <= aes_key_r[APB_DATA_WIDTH-1 : 0];
                                            if(delay_reg1 == 1)
                                            begin
                                                aes_key_r <= aes_key_r >> APB_DATA_WIDTH;
                                            end
                                            en_transfer_r <= 1;
                                        end 
                                    else if( (count == 5'b00011) && (state == SETUP))
                                        begin
                                            en_transfer_r <= 1'b0;
                                            aes_decrypt_write_state <= WRITE_AES_DECRYPT_DATA_IN;                                
                                        end                                                        
                                end
                                
                                WRITE_AES_DECRYPT_DATA_IN:
                                begin
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b01000) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + count*4;
                                            pwdata_r <= aes_text_in_r[APB_DATA_WIDTH-1 : 0];
                                            aes_text_in_r <= aes_text_in_r >> APB_DATA_WIDTH;
                                            en_transfer_r <= 1'b1;
                                        end 
                                    else if( (count == 5'b00111) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 1'b0;
                                            aes_decrypt_write_state <= WRITE_AES_DECRYPT_LOAD;                                
                                        end                                                        
                                end
                                
                                WRITE_AES_DECRYPT_LOAD:
                                begin
                                    pstrb_r <= 4'b0000;
                                    
                                    if( (count < 5'b01001) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + count*4;
                                            pwdata_r <= 32'h00000001;
                                            en_transfer_r <= 1'b1;
                                        end 
                                        
                                    else if( (count == 5'b01001) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + (count - 5'h01)*4;
                                            pwdata_r <= 32'h00000000;
                                            en_transfer_r <= 1'b1;
                                        end
                                        
                                    else if( (count == 5'b01001) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 1'b0;
                                            aes_decrypt_write_state <= WRITE_AES_DECRYPT_K_LOAD;                                    
                                        end 
                                                                                            
                                end
                                
                                WRITE_AES_DECRYPT_K_LOAD:
                                begin
                                    pstrb_r <= 4'b0000;
                                    
                                    if( (count < 5'b01011) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + (count-5'h02)*4;
                                            pwdata_r <= 32'h00010000;
                                            en_transfer_r <= 1'b1;
                                        end 
                                        
                                    else if( (count == 5'b01011) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_WRITE_00 + (count - 5'h03)*4;
                                            pwdata_r <= 32'h00000000;
                                            en_transfer_r <= 1'b1;
                                        end
                                        
                                    else if( (count == 5'b01011) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 1'b0;
//                                            pselx_r <= 0;
                                            operation_complete_r <= 1;
                                        end
                                    
                                    else if( (count == 5'b01011) && (PREADY == 1'b1) )
                                        begin
                                            pselx_r <= 0;
                                        end
                                        
                                    else if( (count == 5'b01100) && (PREADY == 1'b1) )
                                        begin
                                            write_complete_r <= 1;
                                            aes_decrypt_write_state <= WRITE_AES_DECRYPT_INIT;                                    
                                        end 
                                                                                            
                                end
                                
                                default:
                                begin
                                    aes_decrypt_write_state <= WRITE_AES_DECRYPT_INIT;
                                end                        
                              
                            endcase   
                        end
                        
                    AES_DECRYPT_READ: 
                        begin
                            case(aes_decrypt_read_state)
                                
                                READ_AES_DECRYPT_INIT:
                                begin
                                    if( (PREADY == 1) && (slave_sel != 0) )
                                        aes_decrypt_read_state <= READ_AES_DECRYPT_DATA;
                                    en_transfer_r <= 0;
                                end
                                
                                READ_AES_DECRYPT_DATA:
                                begin
                                    pselx_r <= slave_sel;
                                    pwrite_r <= 1'b0;
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b00100) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= (BASE_ADDR_READ_00 + 4*4) + count*4;
                                            decrypt_output_data_r <= {PRDATA, decrypt_output_data_r[AES_INV_CIPH_OUT_WIDTH-1 : APB_DATA_WIDTH]};
                                            en_transfer_r <= 1'b1;
                                        end
                                    else if( (count == 5'b00011) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 0;
//                                            pselx_r <= 0;
                                        end
                                    
                                    else if( (count == 5'b00100) && (PREADY == 1'b1) )
                                            begin
                                                decrypt_output_data_r <= {PRDATA, decrypt_output_data_r[AES_INV_CIPH_OUT_WIDTH-1 : APB_DATA_WIDTH]};
                                                aes_decrypt_read_state <= READ_AES_DECRYPT_DONE;   
                                            end
                                end
                                READ_AES_DECRYPT_DONE:
                                begin
                                    pselx <= 0;
                                    operation_complete_r <= 1;
                                    data_input_ready_r <= 1;
                                    aes_decrypt_read_state <= READ_AES_DECRYPT_INIT;
                                end
                            
                            endcase
                        
                        end 
 //#################################### HASH #################################################  
                    HASH_WRITE:
                        begin
                                pselx_r <= slave_sel;
                                pwrite_r <= 1'b1;
                                case(hash_write_state)
                                    
                                    WRITE_HASH_INIT:
                                    begin
                                        hash_in_r <= hash_in;
                                        if( (PREADY == 1'b1) && (slave_sel != 0) && (write_complete != 1) )
                                            hash_write_state <= WRITE_HASH_DATA_IN;
                                          
                                    end
                                    
                                    WRITE_HASH_DATA_IN:
                                    begin
                                        pstrb_r <= 4'b0000;
                                        if( (count < 5'b10000) && (PREADY == 1'b1) )
                                            begin
                                                paddr_r <= BASE_ADDR_WRITE_01 + count*4;
                                                pwdata_r <= hash_in_r[APB_DATA_WIDTH-1 : 0];
                                                if(delay_reg1 == 1)
                                                begin
                                                    hash_in_r <= hash_in_r >> APB_DATA_WIDTH;
                                                end
                                                en_transfer_r <= 1;
                                            end 
                                        else if( (count == 5'b01111) && (state == SETUP))
                                            begin
                                                en_transfer_r <= 1'b0;
                                                hash_write_state <= WRITE_HASH_GO;                                
                                            end                                                        
                                    end
                                    
                                    WRITE_HASH_GO:
                                    begin
                                        pstrb_r <= 4'b0000;
                                        
                                        if( (count < 5'b10001) && (PREADY == 1'b1) )
                                            begin
                                                paddr_r <= BASE_ADDR_WRITE_01 + count*4;
                                                pwdata_r <= 32'h00000001;
                                                en_transfer_r <= 1'b1;
                                            end 
                                            
                                        else if( (count == 5'b10001) && (PREADY == 1'b1) )
                                            begin
                                                paddr_r <= BASE_ADDR_WRITE_01 + (count - 5'h01)*4;
                                                pwdata_r <= 32'h00000000;
                                                en_transfer_r <= 1'b1;
                                            end
                                            
                                        else if( (count == 5'b10001) && (state == SETUP) )
                                            begin
                                                en_transfer_r <= 1'b0;                                
                                            end
                                            
                                        else if( (count == 5'b10001) && (state == ACCESS) )
                                            begin
//                                                pselx_r <= 0;
                                                operation_complete_r <= 1;                                
                                            end
                                            
                                       else if( (count == 5'b10001) && (PREADY == 1'b1) )
                                            begin
                                                pselx_r <= 0;                               
                                            end
                                            
                                        else if( (count == 5'b10010) && (PREADY == 1'b1) )
                                            begin
                                                write_complete_r <= 1;
                                                hash_write_state <= WRITE_HASH_INIT;                                   
                                            end 
                                                                                                
                                    end
                                    
                                    default:
                                    begin
                                        hash_write_state <= WRITE_HASH_INIT;
                                    end                        
                                  
                                endcase   
                            end

                    HASH_READ: 
                        begin
                            case(hash_read_state)
                                
                                READ_HASH_INIT:
                                begin
                                    if( (PREADY == 1) && (slave_sel != 0) )
                                        hash_read_state <= READ_HASH_DATA;
                                    en_transfer_r <= 0;
                                end
                                
                                READ_HASH_DATA:
                                begin
                                    pselx_r <= slave_sel;
                                    pwrite_r <= 1'b0;
                                    pstrb_r <= 4'b0000;
                                    if( (count < 5'b01000) && (PREADY == 1'b1) )
                                        begin
                                            paddr_r <= BASE_ADDR_READ_01 + count*4;
                                            hash_output_r <= {PRDATA, hash_output_r[HASH_OUT_WIDTH-1 : APB_DATA_WIDTH]};
                                            en_transfer_r <= 1'b1;
                                        end
                                    else if( (count == 5'b00111) && (state == SETUP) )
                                        begin
                                            en_transfer_r <= 0;
//                                            pselx_r <= 0;
                                        end
                                    
                                    else if( (count == 5'b01000) && (PREADY == 1'b1) )
                                            begin
                                                hash_output_r <= {PRDATA, hash_output_r[HASH_OUT_WIDTH-1 : APB_DATA_WIDTH]};
                                                hash_read_state <= READ_HASH_DONE;   
                                            end
                                end
                                
                                READ_HASH_DONE:
                                begin
                                    pselx_r <= 0;
                                    operation_complete_r <= 1;
                                    data_input_ready_r <= 1;
                                    hash_read_state <= READ_HASH_INIT;
                                end
                                
                                default:
                                begin
                                    hash_read_state <= READ_HASH_INIT;
                                end
                            
                            endcase
                        
                        end   
                                   
                endcase
            end

        else if(init_transaction == 0)
            en_transfer_r <= 0;    
            
    end
    
    
    
    
    // APB4 FSM
    always@(posedge PCLK or negedge PRESETn)
    begin
        if( PRESETn == 1'b0 )
            state <= INIT;
        else
            state <= next_state;
    end
    
    always@(*)
    begin
    
        next_state = state;
        paddr = 0;
        pprot = 0;
        pselx = 0;
        pwdata = 0;
        penable = 0;
        pstrb = 0;
        pwrite = 0;
                
        case(state)
            
            INIT:
            begin
                if(en_transfer == 1'b1) begin
                    next_state = IDLE;
                    pselx = pselx_r;
                end
            end
            IDLE:
            begin
                if(en_transfer == 1'b1)
                begin
                    paddr = paddr_r;
                    pprot = pprot_r;
                    pselx = pselx_r;
                    pwrite = pwrite_r;
                    if( pwrite_r == 1'b1 )
                        begin
                            pwdata = pwdata_r;
                            pstrb = pstrb_r;
                        end
                    next_state = SETUP;
                end
            end
            
            SETUP:
            begin
                if(en_transfer == 1'b1)
                begin
                    paddr = paddr_r;
                    pprot = pprot_r;
                    pselx = pselx_r;
                    pwrite = pwrite_r;
                    if( pwrite_r == 1'b1 )
                        begin
                            pwdata = pwdata_r;
                            pstrb = pstrb_r;
                        end
                    penable = 1;
                    next_state = ACCESS;
                end
//                else    
//                    next_state <= IDLE;
                next_state = ACCESS;
            end
            
            ACCESS:
            begin
                paddr = paddr_r;
                pprot = pprot_r;
                pselx = pselx_r;
                pwrite = pwrite_r;
                if( pwrite_r == 1'b1 )
                    begin
                        pwdata = pwdata_r;
                        pstrb = pstrb_r;
                    end
                if( PREADY != 1'b1 )
                    begin
                        penable = 1;
                    end
                else if( PREADY == 1'b1 )
                    begin
                        penable = 0;
                        if( en_transfer == 1'b1 )
                            begin
                                next_state = SETUP;
                            end
                        else
                            begin
                                next_state = INIT; 
                            end
                    end
            end
            
            default:
            begin
                //do nothing 
            end
                        
        endcase
    end
    
    master U_M(
                    .clk(PCLK), 
                    .rstn(PRESETn), 
                    .host_instruction(host_instruction), 
                    .host_data(host_data), 
                    .write_complete(write_complete), 
                    .text_out(aes_text_in), 
                    .key_out(aes_key), 
                    .operation_type(operation_type), 
                    .hash_out(hash_in), 
                    .encrypt_output_data_port(encrypt_output_data), 
                    .decrypt_output_data_port(decrypt_output_data), 
                    .hash_output_port(hash_output), 
                    .data_input_ready(data_input_ready), 
                    .init_transaction(init_transaction), 
                    .start(start), 
                    .operation_done(operation_done),
					.out(out)
					);                   
    
endmodule
